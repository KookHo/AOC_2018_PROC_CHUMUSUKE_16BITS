LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PC IS
PORT
(
		--ativo : IN STD_LOGIC;
		clk :  IN  STD_LOGIC;
		pin :  IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		pout : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
		
	);
END PC;

ARCHITECTURE behavior OF PC IS
BEGIN
	PROCESS(clk)
		BEGIN
			IF rising_edge(clk) THEN
				pout <= pin;
			END IF;
	END PROCESS;
END behavior;